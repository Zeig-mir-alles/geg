`ifndef OVERFLOW_SVH
`define OVERFLOW_SVH

`define FLAGS_OVERFLOW 0

`endif
