`include "execute.svh"

module execute(clk, operation);

input logic clk;
input operation_t operation;

always @(posedge clk) begin

end

endmodule
