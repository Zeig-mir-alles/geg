module registers;

reg [4:0] gprs[31:0];
reg [31:0] flags;
reg [31:0] pc;

endmodule
