`ifndef CACHE_SVH_
`define CACHE_SVH_

`define MEM_OPERATION_READ 0
`define MEM_OPERATION_WRITE 1

`endif
