`include "decode.svh"

module fetch(clk, instruction);
	input logic clk;
	output instruction_t instruction;

	always @(posedge clk) begin

	end
endmodule
